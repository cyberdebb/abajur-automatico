--
-- Curso de FPGA WR Kits Channel
--
--
-- Utilizando o Display de 7 Segmentos
--
--  Truth Table:
--
--                 Entradas    | Saída (segmentos)                                                          
--               D3 D2 D1 D0   |  h g f e d c b a                                                       
--                0  0  0  0   |  0 0 1 1 1 1 1 1                                              
--                0  0  0  1   |  0 0 0 0 0 1 1 0                                                            
--                0  0  1  0   |  0 1 0 1 1 0 1 1                                                             
--                0  0  1  1   |  0 1 0 0 1 1 1 1                                                                   
--                0  1  0  0   |  0 1 1 0 0 1 1 0                                                                           
--                0  1  0  1   |  0 1 1 0 1 1 0 1                                                                              
--                0  1  1  0   |  0 1 1 1 1 1 0 1                                                                             
--                0  1  1  1   |  0 0 0 0 0 1 1 1                                                                                  
--                1  0  0  0   |  0 1 1 1 1 1 1 1                                                       
--                1  0  0  1   |  0 1 1 0 1 1 1 1                                                             
--                                                                                                                        
--


	library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_arith.all;
	use ieee.std_logic_unsigned.all;
	
	
	entity disp7seg is
	port(
	    Data_In          :   in  std_logic_vector(3 downto 0);
        a,b,c,d,e,f,g,h  :  out  std_logic);
		  
   end disp7seg;
	
	
	architecture hardware of disp7seg is
	begin
		process(Data_In)
		begin
		  case Data_In is
-- Applying a low logic level to a segment causes it to light up, and applying a high logic level turns it off.
			when "0000" => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '1'; h <= '1';  -- 0
			when "0001" => a <= '1'; b <= '0'; c <= '0' ; d <= '1'; e <= '1'; f <= '1'; g <= '1'; h <= '1';  -- 1
			when "0010" => a <= '0'; b <= '0'; c <= '1' ; d <= '0'; e <= '0'; f <= '1'; g <= '0'; h <= '1';  -- 2
			when "0011" => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '1'; f <= '1'; g <= '0'; h <= '1';  -- 3 
			when "0100" => a <= '1'; b <= '0'; c <= '0' ; d <= '1'; e <= '1'; f <= '0'; g <= '0'; h <= '1';  -- 4
			when "0101" => a <= '0'; b <= '1'; c <= '0' ; d <= '0'; e <= '1'; f <= '0'; g <= '0'; h <= '1';  -- 5
			when "0110" => a <= '0'; b <= '1'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '1';  -- 6
			when "0111" => a <= '0'; b <= '0'; c <= '0' ; d <= '1'; e <= '1'; f <= '1'; g <= '1'; h <= '1';  -- 7
			when "1000" => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '1';  -- 8
			when "1001" => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '1'; f <= '0'; g <= '0'; h <= '1';  -- 9
			when "1010" => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '0';  -- A
			when "1011" => a <= '1'; b <= '1'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '1';  -- B
			when "1100" => a <= '0'; b <= '1'; c <= '1' ; d <= '0'; e <= '0'; f <= '0'; g <= '1'; h <= '1';  -- C
			when "1101" => a <= '1'; b <= '0'; c <= '0' ; d <= '0'; e <= '0'; f <= '1'; g <= '0'; h <= '1';  -- D
			when "1110" => a <= '1'; b <= '1'; c <= '1' ; d <= '1'; e <= '1'; f <= '1'; g <= '0'; h <= '1';  -- -
			when "1111" => a <= '0'; b <= '1'; c <= '1' ; d <= '1'; e <= '0'; f <= '0'; g <= '0'; h <= '1';  -- F
			when others => a <= '0'; b <= '0'; c <= '0' ; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '0';  -- 
			-- when "0000"   => a <= '1'; b <= '1'; c <= '1'; d <= '1'; e <= '1'; f <= '1'; g <= '0'; h <= '0';
	      	-- when "0001"   => a <= '0'; b <= '1'; c <= '1'; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '0';
			-- when "0010"   => a <= '1'; b <= '1'; c <= '0'; d <= '1'; e <= '1'; f <= '0'; g <= '1'; h <= '0';	
	      	-- when "0011"   => a <= '1'; b <= '1'; c <= '1'; d <= '1'; e <= '0'; f <= '0'; g <= '1'; h <= '0'; 
	      	-- when "0100"   => a <= '0'; b <= '1'; c <= '1'; d <= '0'; e <= '0'; f <= '1'; g <= '1'; h <= '0';	
	      	-- when "0101"   => a <= '1'; b <= '0'; c <= '1'; d <= '1'; e <= '0'; f <= '1'; g <= '1'; h <= '0';	
	      	-- when "0110"   => a <= '1'; b <= '0'; c <= '1'; d <= '1'; e <= '1'; f <= '1'; g <= '1'; h <= '0';	
	      	-- when "0111"   => a <= '1'; b <= '1'; c <= '1'; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '0';	
	      	-- when "1000"   => a <= '1'; b <= '1'; c <= '1'; d <= '1'; e <= '1'; f <= '1'; g <= '1'; h <= '0';
	      	-- when "1001"   => a <= '1'; b <= '1'; c <= '1'; d <= '1'; e <= '0'; f <= '1'; g <= '1'; h <= '0';
			-- when "1110"	  => a <= '1'; b <= '1'; c <= '1'; d <= '1'; e <= '1'; f <= '1'; g <= '0'; h <= '1';		
	      	-- when others   => a <= '0'; b <= '0'; c <= '0'; d <= '0'; e <= '0'; f <= '0'; g <= '0'; h <= '0';	
		end case;
	end process;
		
		
end hardware;
	